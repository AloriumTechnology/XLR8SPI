// *****************************************************
// AVR address constants (localparams)
//  for registers used by Xcelerator Blocks (XBs) 
// *****************************************************

localparam SPCR1_ADDR = 8'hAC;
localparam SPSR1_ADDR = 8'hAD;
localparam SPDR1_ADDR = 8'hAE;

localparam SPCR2_ADDR = 8'hF1;
localparam SPSR2_ADDR = 8'hF2;
localparam SPDR2_ADDR = 8'hF3;
